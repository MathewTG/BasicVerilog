// Simple AND
//----------------------------------
// FileName : simpleand.v
// Type : module
// Author : Mathew T G
// Contact : mathewtg.mec@gmail.com
//------------------
// Date : 15/10/2018
//------------------
// Notes :- Too Simple for a note na ?
//

module simple_and (f,x,y);
input x,y;
output f;
assign f=x&y;
endmodule
